module ALU(
    input wire ALU_control[1:0]
);



endmodule